`ifndef GUARD_GLOBALS
`define GUARD_GLOBALS

`define DATA_W 32
`define OPER_W 32

`endif
